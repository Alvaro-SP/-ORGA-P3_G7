CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
170 0 8 80 10
176 83 1022 713
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
48 C:\Program Files\CircuitMaker 2000 Trial\BOM.DAT
0 7
0 4 0.500000 0.500000
344 179 457 276
42991634 0
0
6 Title:
5 Name:
0
0
0
20
7 Ground~
168 224 424 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7177 0 0
2
5.89311e-315 0
0
14 Logic Display~
6 969 43 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5910 0 0
2
5.89311e-315 0
0
14 Logic Display~
6 951 43 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4350 0 0
2
5.89311e-315 0
0
14 Logic Display~
6 934 43 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3764 0 0
2
5.89311e-315 0
0
14 Logic Display~
6 916 44 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3166 0 0
2
5.89311e-315 0
0
5 7415~
219 676 595 0 4 22
0 8 4 3 9
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U8A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 8 0
1 U
3978 0 0
2
5.89311e-315 0
0
8 2-In OR~
219 738 542 0 3 22
0 10 9 7
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U7C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
9736 0 0
2
5.89311e-315 0
0
9 2-In AND~
219 564 533 0 3 22
0 11 5 10
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
7319 0 0
2
5.89311e-315 0
0
8 2-In OR~
219 493 524 0 3 22
0 13 12 11
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U7B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
6814 0 0
2
5.89311e-315 0
0
8 2-In OR~
219 863 218 0 3 22
0 17 16 14
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U7A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
5585 0 0
2
5.89311e-315 0
0
9 4-In AND~
219 818 260 0 5 22
0 5 4 3 15 16
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U3A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 4 0
1 U
9317 0 0
2
5.89311e-315 0
0
8 3-In OR~
219 668 147 0 4 22
0 12 13 8 18
0
0 0 624 270
4 4075
-14 -24 14 -16
3 U6A
28 -7 49 1
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 6 0
1 U
317 0 0
2
5.89311e-315 0
0
9 2-In AND~
219 755 209 0 3 22
0 18 6 17
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
6624 0 0
2
5.89311e-315 0
0
9 2-In XOR~
219 353 332 0 3 22
0 3 4 19
0
0 0 624 0
5 74F86
-18 -24 17 -16
3 U2A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
6140 0 0
2
5.89311e-315 0
0
7 Ground~
168 373 226 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9118 0 0
2
5.89311e-315 0
0
5 4013~
219 702 361 0 6 22
0 2 14 20 2 15 6
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U1D
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 0 2 2 2 0
1 U
8761 0 0
2
5.89311e-315 0
0
5 4013~
219 566 364 0 6 22
0 2 7 20 2 8 5
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U1C
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 0 2 1 2 0
1 U
3420 0 0
2
5.89311e-315 0
0
5 4013~
219 418 368 0 6 22
0 2 19 20 2 12 4
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U5B
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 0 2 2 1 0
1 U
4545 0 0
2
5.89311e-315 0
0
5 4013~
219 252 369 0 6 22
0 2 13 20 2 13 3
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U5A
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 0 2 1 1 0
1 U
545 0 0
2
5.89311e-315 0
0
7 Pulser~
4 96 352 0 10 12
0 21 22 23 20 0 0 10 10 2
7
0
0 0 4656 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
7476 0 0
2
5.89311e-315 0
0
42
1 0 2 0 0 8192 0 1 0 0 41 3
224 418
224 415
252 415
1 0 3 0 0 8320 0 2 0 0 17 4
969 61
969 71
327 71
327 265
1 0 4 0 0 8320 0 3 0 0 18 4
951 61
951 80
466 80
466 256
1 0 5 0 0 8320 0 4 0 0 19 4
934 61
934 95
615 95
615 247
1 0 6 0 0 4224 0 5 0 0 26 3
916 62
916 296
747 296
3 2 7 0 0 12416 0 7 17 0 0 8
771 542
818 542
818 617
423 617
423 463
511 463
511 328
542 328
3 0 3 0 0 0 0 6 0 0 29 3
652 604
314 604
314 323
2 0 4 0 0 0 0 6 0 0 28 3
652 595
466 595
466 498
1 0 8 0 0 8320 0 6 0 0 25 3
652 586
643 586
643 344
4 2 9 0 0 8320 0 6 7 0 0 4
697 595
708 595
708 551
725 551
3 1 10 0 0 4224 0 8 7 0 0 2
585 533
725 533
2 0 5 0 0 0 0 8 0 0 19 5
540 542
524 542
524 563
615 563
615 327
1 3 11 0 0 4224 0 8 9 0 0 2
540 524
526 524
2 0 12 0 0 8192 0 9 0 0 23 3
480 533
456 533
456 350
1 0 13 0 0 4096 0 9 0 0 31 3
480 515
299 515
299 351
3 2 14 0 0 8336 0 10 16 0 0 6
896 218
902 218
902 456
671 456
671 325
678 325
3 0 3 0 0 0 0 11 0 0 29 3
794 265
326 265
326 323
2 0 4 0 0 0 0 11 0 0 28 3
794 256
466 256
466 332
1 6 5 0 0 0 0 11 17 0 0 4
794 247
615 247
615 328
590 328
4 5 15 0 0 8320 0 11 16 0 0 4
794 274
787 274
787 343
732 343
5 2 16 0 0 8320 0 11 10 0 0 4
839 260
840 260
840 227
850 227
1 3 17 0 0 4224 0 10 13 0 0 2
850 209
776 209
1 5 12 0 0 12416 0 12 18 0 0 5
680 131
680 87
486 87
486 350
448 350
2 0 13 0 0 8320 0 12 0 0 31 5
671 132
671 64
300 64
300 241
299 241
3 5 8 0 0 0 0 12 17 0 0 5
662 131
662 116
643 116
643 346
596 346
2 6 6 0 0 0 0 13 16 0 0 6
731 218
672 218
672 240
747 240
747 325
726 325
4 1 18 0 0 8320 0 12 13 0 0 3
671 177
671 200
731 200
2 6 4 0 0 0 0 14 18 0 0 6
337 341
323 341
323 498
466 498
466 332
442 332
1 6 3 0 0 0 0 14 19 0 0 4
337 323
288 323
288 333
276 333
3 2 19 0 0 4224 0 14 18 0 0 2
386 332
394 332
2 5 13 0 0 0 0 19 19 0 0 6
228 333
213 333
213 241
299 241
299 351
282 351
1 0 2 0 0 12288 0 15 0 0 33 4
373 220
373 209
418 209
418 271
1 0 2 0 0 0 0 18 0 0 35 2
418 311
418 271
1 0 2 0 0 0 0 17 0 0 35 2
566 307
566 271
1 1 2 0 0 8320 0 19 16 0 0 4
252 312
252 271
702 271
702 304
3 0 20 0 0 12288 0 16 0 0 37 4
678 343
659 343
659 442
529 442
3 0 20 0 0 12288 0 17 0 0 38 4
542 346
529 346
529 442
362 442
3 0 20 0 0 12416 0 18 0 0 42 5
394 350
362 350
362 442
164 442
164 351
4 0 2 0 0 0 0 18 0 0 41 2
418 374
418 416
4 0 2 0 0 0 0 17 0 0 41 2
566 370
566 416
4 4 2 0 0 0 0 19 16 0 0 4
252 375
252 416
702 416
702 367
4 3 20 0 0 0 0 20 19 0 0 4
126 352
164 352
164 351
228 351
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
